`define TLAST_PRESENT
`define TSTRB_PRESENT
`define TID_PRESENT
