`include "defines.svh"

module axi_ram 
#(
    parameter ID_W_WIDTH = 4,
    parameter ID_R_WIDTH = 4,
    parameter ADDR_WIDTH = 16,

    parameter AXI_DATA_WIDTH = 32
    `ifdef TID_PRESENT
    ,
    parameter ID_WIDTH = 4
    `endif
    `ifdef TDEST_PRESENT
    ,
    parameter DEST_WIDTH = 4
    `endif
    `ifdef TUSER_PRESENT
    ,
    parameter USER_WIDTH = 4
    `endif,

    parameter BYTE_WIDTH = 8
) (
	input logic clk_i, rst_n_i,
    
    input  axi_mosi_t in_mosi_i,
    output axi_miso_t in_miso_o

);

    `include "axi_type.svh"

    localparam WSRTB_W = AXI_DATA_WIDTH/BYTE_WIDTH;
    
    logic [ADDR_WIDTH-1:0] waddr, raddr;
    logic [BYTE_WIDTH*WSRTB_W-1:0] wdata;
    logic [WSRTB_W-1:0] be;
    logic [BYTE_WIDTH*WSRTB_W-1:0] rdata;

    axi2ram #(
        .ID_W_WIDTH(ID_W_WIDTH),
        .ID_R_WIDTH(ID_R_WIDTH),
        .ADDR_WIDTH(ADDR_WIDTH),

        .AXI_DATA_WIDTH(AXI_DATA_WIDTH)
        `ifdef TID_PRESENT
         ,
        .ID_WIDTH(ID_WIDTH)
        `endif
        `ifdef TDEST_PRESENT
         ,
        .DEST_WIDTH(DEST_WIDTH)
        `endif
        `ifdef TUSER_PRESENT
         ,
        .USER_WIDTH(USER_WIDTH)
        `endif
    
    ) axi (
        .clk_i(clk_i), .rst_n_i(rst_n_i),
        
        .waddr(waddr),
        .raddr(raddr),
        .wdata(wdata),
        .be(be),
        .rdata(rdata),

        .in_mosi_i(in_mosi_i),
        .in_miso_o(in_miso_o)

    );

    generate
        genvar i;
        for (i = 0; i < WSRTB_W; i++) begin : generate_rams
            ram #(
                .ADDR_WIDTH(ADDR_WIDTH),
                .BYTE_WIDTH(BYTE_WIDTH)
            ) coupled_ram (
                .clk_i(clk_i),
                
                .waddr(waddr),
                .raddr(raddr),
                .wdata(wdata[i*BYTE_WIDTH +: BYTE_WIDTH]),
                .we(we & be[i]),
                .rdata(rdata[i*BYTE_WIDTH +: BYTE_WIDTH])

            );
        end
    endgenerate
  
endmodule : axi_ram