`ifndef _DEFINES_
`define _DEFINES_

`define TLAST_PRESENT
`define TSTRB_PRESENT
`define TID_PRESENT

`endif
