`ifndef AXI_TYPE_TEST_SVH
`define AXI_TYPE_TEST_SVH

`include "defines.svh"

parameter ADDR_WIDTH = 16;
parameter ID_R_WIDTH = 4;
parameter ID_W_WIDTH = 4;

`include "axi_type.svh"

`endif
