`define TEST

parameter DATA_WIDTH = 32;

`include "axi_type_test.svh"
`include "axis_type_test.svh"
